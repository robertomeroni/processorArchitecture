`include "constants.v"
`include "dataMemory.v"
`include "dCache.v"

module memoryStage (
		    input clk, rst,
		    input [`WORD_SIZE-1:0] ALUResultM, WriteDataM, PCPlus4M,
		    input [4:0] RdM,
		    // Control ports.
		    input RegWriteM, MemWriteM,
		    input [1:0] ResultSrcM,
		    input ByteAddressM,
		    input ReadEnableM, 

		    // hazard output
		    output [4:0] RdMH,
		    output [0:0] RegWriteMH,
		    output [`WORD_SIZE-1:0] ALUResultW, ReadDataW, PCPlus4W,
		    output [4:0] RdW,
		    output RegWriteW,
		    output [1:0] ResultSrcW,
		    output CacheStall
		    );

   // Internal wires and registers.
   wire [`WORD_SIZE-1:0] ReadDataM;
   wire Ready;
   wire [`CACHE_LINE_SIZE-1:0] MemLine;
   wire MemRead;
   wire CacheStall;
   wire [`WORD_SIZE-1:0] AMem;


   reg [`WORD_SIZE-1:0] ALUResultM_reg, ReadDataM_reg, PCPlus4M_reg;
   reg [4:0] RdM_reg;

   // Control signals and registers.
   reg RegWriteM_reg;
   reg [1:0] ResultSrcM_reg;

   // Modules.
   dataMemory Data_Memory (
			   .clk(clk),
			   .rst(rst),
			   .WE(MemWriteM),
			   .WD(WriteDataM),
			   .A(ALUResultM),
			   .ByteAddress(ByteAddressM),
			   .Ready(Ready),
			   .Line(MemLine),
			   .Read(MemRead)
			   );

   dCache Data_Cache (
		      .clk(clk),
		      .rst(rst),
		      .A(ALUResultM),
		      .ReadEnable(ReadEnableM),
		      .AMem(AMem),
		      .MemLine(MemLine),
		      .MemReady(Ready),
		      .MemRead(MemRead),
		      .Value(ReadDataM),
		      .CacheStall(CacheStall)
		      );

   // Behavior.
   // TODO: make memory access take 5 clocks as per the project statement
   always @(posedge clk or posedge rst) begin
      if (rst) begin
         ALUResultM_reg <= 0;
         ReadDataM_reg <= 0;
         PCPlus4M_reg <= 0;
         RdM_reg <= 0;
         RegWriteM_reg <= 0;
         ResultSrcM_reg <= 0;
      end else begin
         ALUResultM_reg <= ALUResultM;
         ReadDataM_reg <= ReadDataM;
         PCPlus4M_reg <= PCPlus4M;
         RdM_reg <= RdM;
         RegWriteM_reg <= RegWriteM;
         ResultSrcM_reg <= ResultSrcM;
      end
      #4;
      $display("--- MEMORY STAGE ---");
      $display("MemWriteM = %1b", MemWriteM);
      $display("ALUResultM = %32b", ALUResultM);
      $display("RegWriteM = %1b", RegWriteM);
      $display("--- ------ ----- ---");
      $display("ReadDataW = %32b", ReadDataW);
   end

   // Outputs.
   assign RdMH = RdM;
   assign RegWriteMH = RegWriteM;
   assign ALUResultW = ALUResultM_reg;
   assign ReadDataW = ReadDataM_reg;
   assign PCPlus4W = PCPlus4M_reg;
   assign RdW = RdM_reg;
   assign RegWriteW = RegWriteM_reg;
   assign ResultSrcW = ResultSrcM_reg;
endmodule

