`include "constants.v"

module controlUnit (
    input [6:0] Op,
    input [2:0] funct3,
    input funct7,
    output RegWrite, MemWrite, Jump, Branch, ALUSrc,
    output [1:0] ResultSrc, ImmSrc,
    output [2:0] ALUControl
);

// TODO: Complete this module.
    
)