`include "constants.v"

module controlUnit (
    input [6:0] Op,
    input [2:0] funct3,
    input funct7,
    output RegWrite,
    output [1:0] ResultSrc,
    output MemWrite,
    output Jump,
    output Branch,
    output [2:0] ALUControl,
    output ALUSrc,
    output [1:0] ImmSrc,
    );

// TODO: Complete this module.
    
)