`include "constants.v"

module memoryStage(clk, rst, ALUResultM, WriteDataM, RdM, PCPlus4M, RD)